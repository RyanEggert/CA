module hw1test;
initial begin
$display("Hello, CompArch!");
end
endmodule
